-- Synthesisable design for a sine wave generator
-- Copyright Doulos Ltd
-- SD, 07 Aug 2003
library ieee;
use ieee.std_logic_1164.all;

package sine_package is

  constant max_table_value: integer := 255;
  subtype table_value_type is integer range 0 to max_table_value;

  constant max_table_index: integer := 511;
  subtype table_index_type is integer range 0 to max_table_index;

  subtype sine_vector_type is std_logic_vector( 8 downto 0 );

  function get_table_value (table_index: table_index_type) return table_value_type;

end;

package body sine_package is

  function get_table_value (table_index: table_index_type) return table_value_type is
    variable table_value: table_value_type;
  begin
    case table_index is
      when 0 =>
        table_value := 0;
      when 1 =>
        table_value := 1;
      when 2 =>
        table_value := 2;
      when 3 =>
        table_value := 3;
      when 4 =>
        table_value := 4;
      when 5 =>
        table_value := 4;
      when 6 =>
        table_value := 5;
      when 7 =>
        table_value := 6;
      when 8 =>
        table_value := 7;
      when 9 =>
        table_value := 7;
      when 10 =>
        table_value := 8;
      when 11 =>
        table_value := 9;
      when 12 =>
        table_value := 10;
      when 13 =>
        table_value := 11;
      when 14 =>
        table_value := 11;
      when 15 =>
        table_value := 12;
      when 16 =>
        table_value := 13;
      when 17 =>
        table_value := 14;
      when 18 =>
        table_value := 14;
      when 19 =>
        table_value := 15;
      when 20 =>
        table_value := 16;
      when 21 =>
        table_value := 17;
      when 22 =>
        table_value := 18;
      when 23 =>
        table_value := 18;
      when 24 =>
        table_value := 19;
      when 25 =>
        table_value := 20;
      when 26 =>
        table_value := 21;
      when 27 =>
        table_value := 21;
      when 28 =>
        table_value := 22;
      when 29 =>
        table_value := 23;
      when 30 =>
        table_value := 24;
      when 31 =>
        table_value := 25;
      when 32 =>
        table_value := 25;
      when 33 =>
        table_value := 26;
      when 34 =>
        table_value := 27;
      when 35 =>
        table_value := 28;
      when 36 =>
        table_value := 28;
      when 37 =>
        table_value := 29;
      when 38 =>
        table_value := 30;
      when 39 =>
        table_value := 31;
      when 40 =>
        table_value := 32;
      when 41 =>
        table_value := 32;
      when 42 =>
        table_value := 33;
      when 43 =>
        table_value := 34;
      when 44 =>
        table_value := 35;
      when 45 =>
        table_value := 35;
      when 46 =>
        table_value := 36;
      when 47 =>
        table_value := 37;
      when 48 =>
        table_value := 38;
      when 49 =>
        table_value := 39;
      when 50 =>
        table_value := 39;
      when 51 =>
        table_value := 40;
      when 52 =>
        table_value := 41;
      when 53 =>
        table_value := 42;
      when 54 =>
        table_value := 42;
      when 55 =>
        table_value := 43;
      when 56 =>
        table_value := 44;
      when 57 =>
        table_value := 45;
      when 58 =>
        table_value := 46;
      when 59 =>
        table_value := 46;
      when 60 =>
        table_value := 47;
      when 61 =>
        table_value := 48;
      when 62 =>
        table_value := 49;
      when 63 =>
        table_value := 49;
      when 64 =>
        table_value := 50;
      when 65 =>
        table_value := 51;
      when 66 =>
        table_value := 52;
      when 67 =>
        table_value := 52;
      when 68 =>
        table_value := 53;
      when 69 =>
        table_value := 54;
      when 70 =>
        table_value := 55;
      when 71 =>
        table_value := 55;
      when 72 =>
        table_value := 56;
      when 73 =>
        table_value := 57;
      when 74 =>
        table_value := 58;
      when 75 =>
        table_value := 59;
      when 76 =>
        table_value := 59;
      when 77 =>
        table_value := 60;
      when 78 =>
        table_value := 61;
      when 79 =>
        table_value := 62;
      when 80 =>
        table_value := 62;
      when 81 =>
        table_value := 63;
      when 82 =>
        table_value := 64;
      when 83 =>
        table_value := 65;
      when 84 =>
        table_value := 65;
      when 85 =>
        table_value := 66;
      when 86 =>
        table_value := 67;
      when 87 =>
        table_value := 68;
      when 88 =>
        table_value := 68;
      when 89 =>
        table_value := 69;
      when 90 =>
        table_value := 70;
      when 91 =>
        table_value := 71;
      when 92 =>
        table_value := 71;
      when 93 =>
        table_value := 72;
      when 94 =>
        table_value := 73;
      when 95 =>
        table_value := 74;
      when 96 =>
        table_value := 74;
      when 97 =>
        table_value := 75;
      when 98 =>
        table_value := 76;
      when 99 =>
        table_value := 77;
      when 100 =>
        table_value := 77;
      when 101 =>
        table_value := 78;
      when 102 =>
        table_value := 79;
      when 103 =>
        table_value := 80;
      when 104 =>
        table_value := 80;
      when 105 =>
        table_value := 81;
      when 106 =>
        table_value := 82;
      when 107 =>
        table_value := 83;
      when 108 =>
        table_value := 83;
      when 109 =>
        table_value := 84;
      when 110 =>
        table_value := 85;
      when 111 =>
        table_value := 86;
      when 112 =>
        table_value := 86;
      when 113 =>
        table_value := 87;
      when 114 =>
        table_value := 88;
      when 115 =>
        table_value := 88;
      when 116 =>
        table_value := 89;
      when 117 =>
        table_value := 90;
      when 118 =>
        table_value := 91;
      when 119 =>
        table_value := 91;
      when 120 =>
        table_value := 92;
      when 121 =>
        table_value := 93;
      when 122 =>
        table_value := 94;
      when 123 =>
        table_value := 94;
      when 124 =>
        table_value := 95;
      when 125 =>
        table_value := 96;
      when 126 =>
        table_value := 96;
      when 127 =>
        table_value := 97;
      when 128 =>
        table_value := 98;
      when 129 =>
        table_value := 99;
      when 130 =>
        table_value := 99;
      when 131 =>
        table_value := 100;
      when 132 =>
        table_value := 101;
      when 133 =>
        table_value := 102;
      when 134 =>
        table_value := 102;
      when 135 =>
        table_value := 103;
      when 136 =>
        table_value := 104;
      when 137 =>
        table_value := 104;
      when 138 =>
        table_value := 105;
      when 139 =>
        table_value := 106;
      when 140 =>
        table_value := 107;
      when 141 =>
        table_value := 107;
      when 142 =>
        table_value := 108;
      when 143 =>
        table_value := 109;
      when 144 =>
        table_value := 109;
      when 145 =>
        table_value := 110;
      when 146 =>
        table_value := 111;
      when 147 =>
        table_value := 111;
      when 148 =>
        table_value := 112;
      when 149 =>
        table_value := 113;
      when 150 =>
        table_value := 114;
      when 151 =>
        table_value := 114;
      when 152 =>
        table_value := 115;
      when 153 =>
        table_value := 116;
      when 154 =>
        table_value := 116;
      when 155 =>
        table_value := 117;
      when 156 =>
        table_value := 118;
      when 157 =>
        table_value := 118;
      when 158 =>
        table_value := 119;
      when 159 =>
        table_value := 120;
      when 160 =>
        table_value := 121;
      when 161 =>
        table_value := 121;
      when 162 =>
        table_value := 122;
      when 163 =>
        table_value := 123;
      when 164 =>
        table_value := 123;
      when 165 =>
        table_value := 124;
      when 166 =>
        table_value := 125;
      when 167 =>
        table_value := 125;
      when 168 =>
        table_value := 126;
      when 169 =>
        table_value := 127;
      when 170 =>
        table_value := 127;
      when 171 =>
        table_value := 128;
      when 172 =>
        table_value := 129;
      when 173 =>
        table_value := 129;
      when 174 =>
        table_value := 130;
      when 175 =>
        table_value := 131;
      when 176 =>
        table_value := 131;
      when 177 =>
        table_value := 132;
      when 178 =>
        table_value := 133;
      when 179 =>
        table_value := 133;
      when 180 =>
        table_value := 134;
      when 181 =>
        table_value := 135;
      when 182 =>
        table_value := 135;
      when 183 =>
        table_value := 136;
      when 184 =>
        table_value := 137;
      when 185 =>
        table_value := 137;
      when 186 =>
        table_value := 138;
      when 187 =>
        table_value := 139;
      when 188 =>
        table_value := 139;
      when 189 =>
        table_value := 140;
      when 190 =>
        table_value := 141;
      when 191 =>
        table_value := 141;
      when 192 =>
        table_value := 142;
      when 193 =>
        table_value := 143;
      when 194 =>
        table_value := 143;
      when 195 =>
        table_value := 144;
      when 196 =>
        table_value := 145;
      when 197 =>
        table_value := 145;
      when 198 =>
        table_value := 146;
      when 199 =>
        table_value := 147;
      when 200 =>
        table_value := 147;
      when 201 =>
        table_value := 148;
      when 202 =>
        table_value := 148;
      when 203 =>
        table_value := 149;
      when 204 =>
        table_value := 150;
      when 205 =>
        table_value := 150;
      when 206 =>
        table_value := 151;
      when 207 =>
        table_value := 152;
      when 208 =>
        table_value := 152;
      when 209 =>
        table_value := 153;
      when 210 =>
        table_value := 153;
      when 211 =>
        table_value := 154;
      when 212 =>
        table_value := 155;
      when 213 =>
        table_value := 155;
      when 214 =>
        table_value := 156;
      when 215 =>
        table_value := 157;
      when 216 =>
        table_value := 157;
      when 217 =>
        table_value := 158;
      when 218 =>
        table_value := 158;
      when 219 =>
        table_value := 159;
      when 220 =>
        table_value := 160;
      when 221 =>
        table_value := 160;
      when 222 =>
        table_value := 161;
      when 223 =>
        table_value := 161;
      when 224 =>
        table_value := 162;
      when 225 =>
        table_value := 163;
      when 226 =>
        table_value := 163;
      when 227 =>
        table_value := 164;
      when 228 =>
        table_value := 164;
      when 229 =>
        table_value := 165;
      when 230 =>
        table_value := 166;
      when 231 =>
        table_value := 166;
      when 232 =>
        table_value := 167;
      when 233 =>
        table_value := 167;
      when 234 =>
        table_value := 168;
      when 235 =>
        table_value := 169;
      when 236 =>
        table_value := 169;
      when 237 =>
        table_value := 170;
      when 238 =>
        table_value := 170;
      when 239 =>
        table_value := 171;
      when 240 =>
        table_value := 172;
      when 241 =>
        table_value := 172;
      when 242 =>
        table_value := 173;
      when 243 =>
        table_value := 173;
      when 244 =>
        table_value := 174;
      when 245 =>
        table_value := 174;
      when 246 =>
        table_value := 175;
      when 247 =>
        table_value := 176;
      when 248 =>
        table_value := 176;
      when 249 =>
        table_value := 177;
      when 250 =>
        table_value := 177;
      when 251 =>
        table_value := 178;
      when 252 =>
        table_value := 178;
      when 253 =>
        table_value := 179;
      when 254 =>
        table_value := 179;
      when 255 =>
        table_value := 180;
      when 256 =>
        table_value := 181;
      when 257 =>
        table_value := 181;
      when 258 =>
        table_value := 182;
      when 259 =>
        table_value := 182;
      when 260 =>
        table_value := 183;
      when 261 =>
        table_value := 183;
      when 262 =>
        table_value := 184;
      when 263 =>
        table_value := 184;
      when 264 =>
        table_value := 185;
      when 265 =>
        table_value := 185;
      when 266 =>
        table_value := 186;
      when 267 =>
        table_value := 187;
      when 268 =>
        table_value := 187;
      when 269 =>
        table_value := 188;
      when 270 =>
        table_value := 188;
      when 271 =>
        table_value := 189;
      when 272 =>
        table_value := 189;
      when 273 =>
        table_value := 190;
      when 274 =>
        table_value := 190;
      when 275 =>
        table_value := 191;
      when 276 =>
        table_value := 191;
      when 277 =>
        table_value := 192;
      when 278 =>
        table_value := 192;
      when 279 =>
        table_value := 193;
      when 280 =>
        table_value := 193;
      when 281 =>
        table_value := 194;
      when 282 =>
        table_value := 194;
      when 283 =>
        table_value := 195;
      when 284 =>
        table_value := 195;
      when 285 =>
        table_value := 196;
      when 286 =>
        table_value := 196;
      when 287 =>
        table_value := 197;
      when 288 =>
        table_value := 197;
      when 289 =>
        table_value := 198;
      when 290 =>
        table_value := 198;
      when 291 =>
        table_value := 199;
      when 292 =>
        table_value := 199;
      when 293 =>
        table_value := 200;
      when 294 =>
        table_value := 200;
      when 295 =>
        table_value := 201;
      when 296 =>
        table_value := 201;
      when 297 =>
        table_value := 202;
      when 298 =>
        table_value := 202;
      when 299 =>
        table_value := 203;
      when 300 =>
        table_value := 203;
      when 301 =>
        table_value := 204;
      when 302 =>
        table_value := 204;
      when 303 =>
        table_value := 205;
      when 304 =>
        table_value := 205;
      when 305 =>
        table_value := 206;
      when 306 =>
        table_value := 206;
      when 307 =>
        table_value := 206;
      when 308 =>
        table_value := 207;
      when 309 =>
        table_value := 207;
      when 310 =>
        table_value := 208;
      when 311 =>
        table_value := 208;
      when 312 =>
        table_value := 209;
      when 313 =>
        table_value := 209;
      when 314 =>
        table_value := 210;
      when 315 =>
        table_value := 210;
      when 316 =>
        table_value := 210;
      when 317 =>
        table_value := 211;
      when 318 =>
        table_value := 211;
      when 319 =>
        table_value := 212;
      when 320 =>
        table_value := 212;
      when 321 =>
        table_value := 213;
      when 322 =>
        table_value := 213;
      when 323 =>
        table_value := 214;
      when 324 =>
        table_value := 214;
      when 325 =>
        table_value := 214;
      when 326 =>
        table_value := 215;
      when 327 =>
        table_value := 215;
      when 328 =>
        table_value := 216;
      when 329 =>
        table_value := 216;
      when 330 =>
        table_value := 216;
      when 331 =>
        table_value := 217;
      when 332 =>
        table_value := 217;
      when 333 =>
        table_value := 218;
      when 334 =>
        table_value := 218;
      when 335 =>
        table_value := 219;
      when 336 =>
        table_value := 219;
      when 337 =>
        table_value := 219;
      when 338 =>
        table_value := 220;
      when 339 =>
        table_value := 220;
      when 340 =>
        table_value := 221;
      when 341 =>
        table_value := 221;
      when 342 =>
        table_value := 221;
      when 343 =>
        table_value := 222;
      when 344 =>
        table_value := 222;
      when 345 =>
        table_value := 222;
      when 346 =>
        table_value := 223;
      when 347 =>
        table_value := 223;
      when 348 =>
        table_value := 224;
      when 349 =>
        table_value := 224;
      when 350 =>
        table_value := 224;
      when 351 =>
        table_value := 225;
      when 352 =>
        table_value := 225;
      when 353 =>
        table_value := 225;
      when 354 =>
        table_value := 226;
      when 355 =>
        table_value := 226;
      when 356 =>
        table_value := 227;
      when 357 =>
        table_value := 227;
      when 358 =>
        table_value := 227;
      when 359 =>
        table_value := 228;
      when 360 =>
        table_value := 228;
      when 361 =>
        table_value := 228;
      when 362 =>
        table_value := 229;
      when 363 =>
        table_value := 229;
      when 364 =>
        table_value := 229;
      when 365 =>
        table_value := 230;
      when 366 =>
        table_value := 230;
      when 367 =>
        table_value := 230;
      when 368 =>
        table_value := 231;
      when 369 =>
        table_value := 231;
      when 370 =>
        table_value := 231;
      when 371 =>
        table_value := 232;
      when 372 =>
        table_value := 232;
      when 373 =>
        table_value := 232;
      when 374 =>
        table_value := 233;
      when 375 =>
        table_value := 233;
      when 376 =>
        table_value := 233;
      when 377 =>
        table_value := 234;
      when 378 =>
        table_value := 234;
      when 379 =>
        table_value := 234;
      when 380 =>
        table_value := 235;
      when 381 =>
        table_value := 235;
      when 382 =>
        table_value := 235;
      when 383 =>
        table_value := 235;
      when 384 =>
        table_value := 236;
      when 385 =>
        table_value := 236;
      when 386 =>
        table_value := 236;
      when 387 =>
        table_value := 237;
      when 388 =>
        table_value := 237;
      when 389 =>
        table_value := 237;
      when 390 =>
        table_value := 237;
      when 391 =>
        table_value := 238;
      when 392 =>
        table_value := 238;
      when 393 =>
        table_value := 238;
      when 394 =>
        table_value := 239;
      when 395 =>
        table_value := 239;
      when 396 =>
        table_value := 239;
      when 397 =>
        table_value := 239;
      when 398 =>
        table_value := 240;
      when 399 =>
        table_value := 240;
      when 400 =>
        table_value := 240;
      when 401 =>
        table_value := 240;
      when 402 =>
        table_value := 241;
      when 403 =>
        table_value := 241;
      when 404 =>
        table_value := 241;
      when 405 =>
        table_value := 242;
      when 406 =>
        table_value := 242;
      when 407 =>
        table_value := 242;
      when 408 =>
        table_value := 242;
      when 409 =>
        table_value := 242;
      when 410 =>
        table_value := 243;
      when 411 =>
        table_value := 243;
      when 412 =>
        table_value := 243;
      when 413 =>
        table_value := 243;
      when 414 =>
        table_value := 244;
      when 415 =>
        table_value := 244;
      when 416 =>
        table_value := 244;
      when 417 =>
        table_value := 244;
      when 418 =>
        table_value := 245;
      when 419 =>
        table_value := 245;
      when 420 =>
        table_value := 245;
      when 421 =>
        table_value := 245;
      when 422 =>
        table_value := 245;
      when 423 =>
        table_value := 246;
      when 424 =>
        table_value := 246;
      when 425 =>
        table_value := 246;
      when 426 =>
        table_value := 246;
      when 427 =>
        table_value := 246;
      when 428 =>
        table_value := 247;
      when 429 =>
        table_value := 247;
      when 430 =>
        table_value := 247;
      when 431 =>
        table_value := 247;
      when 432 =>
        table_value := 247;
      when 433 =>
        table_value := 248;
      when 434 =>
        table_value := 248;
      when 435 =>
        table_value := 248;
      when 436 =>
        table_value := 248;
      when 437 =>
        table_value := 248;
      when 438 =>
        table_value := 249;
      when 439 =>
        table_value := 249;
      when 440 =>
        table_value := 249;
      when 441 =>
        table_value := 249;
      when 442 =>
        table_value := 249;
      when 443 =>
        table_value := 249;
      when 444 =>
        table_value := 250;
      when 445 =>
        table_value := 250;
      when 446 =>
        table_value := 250;
      when 447 =>
        table_value := 250;
      when 448 =>
        table_value := 250;
      when 449 =>
        table_value := 250;
      when 450 =>
        table_value := 250;
      when 451 =>
        table_value := 251;
      when 452 =>
        table_value := 251;
      when 453 =>
        table_value := 251;
      when 454 =>
        table_value := 251;
      when 455 =>
        table_value := 251;
      when 456 =>
        table_value := 251;
      when 457 =>
        table_value := 251;
      when 458 =>
        table_value := 252;
      when 459 =>
        table_value := 252;
      when 460 =>
        table_value := 252;
      when 461 =>
        table_value := 252;
      when 462 =>
        table_value := 252;
      when 463 =>
        table_value := 252;
      when 464 =>
        table_value := 252;
      when 465 =>
        table_value := 252;
      when 466 =>
        table_value := 253;
      when 467 =>
        table_value := 253;
      when 468 =>
        table_value := 253;
      when 469 =>
        table_value := 253;
      when 470 =>
        table_value := 253;
      when 471 =>
        table_value := 253;
      when 472 =>
        table_value := 253;
      when 473 =>
        table_value := 253;
      when 474 =>
        table_value := 253;
      when 475 =>
        table_value := 253;
      when 476 =>
        table_value := 253;
      when 477 =>
        table_value := 254;
      when 478 =>
        table_value := 254;
      when 479 =>
        table_value := 254;
      when 480 =>
        table_value := 254;
      when 481 =>
        table_value := 254;
      when 482 =>
        table_value := 254;
      when 483 =>
        table_value := 254;
      when 484 =>
        table_value := 254;
      when 485 =>
        table_value := 254;
      when 486 =>
        table_value := 254;
      when 487 =>
        table_value := 254;
      when 488 =>
        table_value := 254;
      when 489 =>
        table_value := 254;
      when 490 =>
        table_value := 254;
      when 491 =>
        table_value := 254;
      when 492 =>
        table_value := 255;
      when 493 =>
        table_value := 255;
      when 494 =>
        table_value := 255;
      when 495 =>
        table_value := 255;
      when 496 =>
        table_value := 255;
      when 497 =>
        table_value := 255;
      when 498 =>
        table_value := 255;
      when 499 =>
        table_value := 255;
      when 500 =>
        table_value := 255;
      when 501 =>
        table_value := 255;
      when 502 =>
        table_value := 255;
      when 503 =>
        table_value := 255;
      when 504 =>
        table_value := 255;
      when 505 =>
        table_value := 255;
      when 506 =>
        table_value := 255;
      when 507 =>
        table_value := 255;
      when 508 =>
        table_value := 255;
      when 509 =>
        table_value := 255;
      when 510 =>
        table_value := 255;
      when 511 =>
        table_value := 255;
    end case;
    return table_value;
  end;

end;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.sine_package.all;

entity sine_wave is
  port( clock, reset, enable: in std_logic;
        wave_out: out sine_vector_type);
end;

architecture arch1 of sine_wave is
  type state_type is ( counting_up, change_down, counting_down, change_up );
  signal state, next_state: state_type;
  signal table_index: table_index_type;
  signal positive_cycle: boolean;
begin

  process( clock, reset )
  begin
    if reset = '1' then
      state <= counting_up;
    elsif rising_edge( clock ) then
      if enable = '1' then
        state <= next_state;
      end if;
    end if;
  end process;

  process( state, table_index )
  begin
    next_state <= state;
    case state is
      when counting_up =>
        if table_index = max_table_index then
          next_state <= change_down;
        end if;
      when change_down =>
        next_state <= counting_down;
      when counting_down =>
        if table_index = 0 then
          next_state <= change_up;
        end if;
      when others => -- change_up
        next_state <= counting_up;
    end case;
  end process;

  process( clock, reset )
  begin
    if reset = '1' then
      table_index <= 0;
      positive_cycle <= true;
    elsif rising_edge( clock ) then
      if enable = '1' then
        case next_state is
          when counting_up =>
            table_index <= table_index + 1;
          when counting_down =>
            table_index <= table_index - 1;
          when change_up =>
            positive_cycle <= not positive_cycle;
          when others =>
            -- nothing to do
        end case;
      end if;
    end if;
  end process;

  process( table_index, positive_cycle )
    variable table_value: table_value_type;
  begin
    table_value := get_table_value( table_index );
    if positive_cycle then
      wave_out <= std_logic_vector(to_signed(table_value,sine_vector_type'length));
    else
      wave_out <= std_logic_vector(to_signed(-table_value,sine_vector_type'length));
    end if;
  end process;

end;
